package svutest_core_pkg;
    interface class protocol;
        pure virtual task run ();
    endclass
endpackage
