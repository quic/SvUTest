// Copyright (c) 2024 Qualcomm Innovation Center, Inc. All rights reserved.
// SPDX-License-Identifier: BSD-3-Clause-Clear

package svutest_core_pkg;
    interface class protocol;
        pure virtual task run ();
    endclass
endpackage
