// Copyright (c) Qualcomm Technologies, Inc. and/or its subsidiaries.
// SPDX-License-Identifier: BSD-3-Clause-Clear

`ifndef SVUTEST_CORE_SVH
`define SVUTEST_CORE_SVH

interface class protocol;
    pure virtual task run ();
endclass

`endif
