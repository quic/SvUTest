// Copyright (c) 2024 Qualcomm Innovation Center, Inc. All rights reserved.
// SPDX-License-Identifier: BSD-3-Clause-Clear

package svutest_pkg;
    `include "svutest_core.svh"
    `include "svutest_injector.svh"
    `include "svutest_extractor.svh"
    `include "svutest_test.svh"
    `include "svutest_testlist.svh"
endpackage
