// Copyright (c) 2024 Qualcomm Innovation Center, Inc. All rights reserved.
// SPDX-License-Identifier: BSD-3-Clause-Clear

`ifndef SVUTEST_CORE_SVH
`define SVUTEST_CORE_SVH

interface class protocol;
    pure virtual task run ();
endclass

`endif
